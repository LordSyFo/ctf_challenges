
module chip ();

wire n1, n2, io_12_31_1, n112, n114, n137, n138, n139, n140, n141;
wire n142, n143, n144, n145, n146, n147, n148, n155, n156, n158;
wire n159, n176, n180, n183, n184, n185, n187, n188, n189, n190;
wire n191, n192, n193, n194, n195, n196, n197, n199, n200, n201;
wire n202, n203, n204, n205, io_16_0_0, n223, n224, n225, n239, n240;
wire n241, n242, n243, n244, n245, io_17_0_0, n275, n276, n277, n278;
wire n279, n280, n281, n282, n283, n284, n285, n286, n287, n288;
wire n289, n290, n291, n292, n293, n294, n295, n296, n297, n298;
wire n299, n300, n301, n302, n303, n304, n305, n306, n307, n308;
wire n309, n310, n311, n312, n313, n314, n315, n316, n317, n318;
wire n319, n320, n321, n322, n323, n324, n325, n326, n327, n328;
wire n329, n330, n331, n332, n333, n334, n335, n336, n337, n338;
wire n339, n340, n341, n342, n343, n344, n345, n346, n347, n348;
wire n349, n350, n351, n352, n353, n354, n355, n356, n357, n358;
wire n359, n360, n361, n362, n363, n364, n365, n366, n367, n368;
wire n369, n370, n371, n372, n373, n374, n375, n376, n377, n378;
wire n379, n380, n381, n382, n383, n384, n385, n386, n387, n388;
wire n389, n390, n391, n392, n393, n394, n395, n396, n397, n398;
wire n399, n400, n401, n402, n403, n404, n405, n406, n407, n408;
wire n409, n410, n411, n412, n413, n414, n415, n416, n417, n418;
wire n419, n420, n421, n422, n423, n424, n425, n426, n427, n428;
wire n429, n430, n431, n432, n433, n434, n435, n436, n437, n438;
wire n439, n440, n441, n442, n443, n444, n445, n446, n447, n448;
wire n449, n450, n451, n452, n453, n454, n455, n456, n457, n458;
wire n459, n460, n461, n462, n463, n464, n465, n466, n467, n468;
wire n469, n470, n471, n472, n473, n474, n475, n476, n477, n478;
wire n479, n480, n481, n482, n483, n484, n485, n486, n487, n488;
wire n489, n490, n491, n492, n493, n494, n495, n496, n497, n498;
wire n499, n500, n501, n502, n503, n504, n505, n506, n507, n508;
wire n509, n510, n511, n512, n513, n514, n515, n516, n517, n518;
wire n519, n520, n521, n522, n523, n524, n525, n526, n527, n528;
wire n529, n530, n531, n532, n533, n534, n535, n536, n537, n538;
wire n539, n540;
reg n4 = 0, n5 = 0, n6 = 0, n7 = 0, n8 = 0, n9 = 0, n10 = 0, n11 = 0, n12 = 0, n13 = 0;
reg n14 = 0, n15 = 0, n16 = 0, n17 = 0, n18 = 0, n19 = 0, n20 = 0, n21 = 0, n22 = 0, n23 = 0;
reg n24 = 0, n25 = 0, n26 = 0, n27 = 0, n28 = 0, n29 = 0, n30 = 0, n31 = 0, n32 = 0, n33 = 0;
reg n34 = 0, n35 = 0, n36 = 0, n37 = 0, n38 = 0, n39 = 0, n40 = 0, n41 = 0, n42 = 0, n43 = 0;
reg n44 = 0, n45 = 0, n46 = 0, n47 = 0, n48 = 0, n49 = 0, n50 = 0, n51 = 0, n52 = 0, n53 = 0;
reg n54 = 0, n55 = 0, n56 = 0, n57 = 0, n58 = 0, n59 = 0, n60 = 0, n61 = 0, n62 = 0, n63 = 0;
reg n64 = 0, n65 = 0, n66 = 0, n67 = 0, n68 = 0, n69 = 0, n70 = 0, n71 = 0, n72 = 0, n73 = 0;
reg n74 = 0, n75 = 0, n76 = 0, n77 = 0, n78 = 0, n79 = 0, n80 = 0, n81 = 0, n82 = 0, n83 = 0;
reg n84 = 0, n85 = 0, n86 = 0, n87 = 0, n88 = 0, n89 = 0, n90 = 0, n91 = 0, n92 = 0, n93 = 0;
reg n94 = 0, n95 = 0, n96 = 0, n97 = 0, n98 = 0, n99 = 0, n100 = 0, n101 = 0, n102 = 0, n103 = 0;
reg n104 = 0, n105 = 0, n106 = 0, n107 = 0, n108 = 0, n109 = 0, n110 = 0, n111 = 0, n113 = 0, n115 = 0;
reg n116 = 0, n117 = 0, n118 = 0, n119 = 0, n120 = 0, n121 = 0, n122 = 0, n123 = 0, n124 = 0, n125 = 0;
reg n126 = 0, n127 = 0, n128 = 0, n129 = 0, n130 = 0, n131 = 0, n132 = 0, n133 = 0, n134 = 0, n135 = 0;
reg n136 = 0, n149 = 0, n150 = 0, n151 = 0, n152 = 0, n153 = 0, n154 = 0, n157 = 0, n160 = 0, n161 = 0;
reg n162 = 0, n163 = 0, n164 = 0, n165 = 0, n166 = 0, n167 = 0, n168 = 0, n169 = 0, n170 = 0, n171 = 0;
reg n172 = 0, n173 = 0, n174 = 0, n175 = 0, n177 = 0, n178 = 0, n179 = 0, n181 = 0, n182 = 0, n186 = 0;
reg n198 = 0, n206 = 0, n208 = 0, n209 = 0, n210 = 0, n211 = 0, n212 = 0, n213 = 0, n214 = 0, n215 = 0;
reg n216 = 0, n217 = 0, n218 = 0, n219 = 0, n220 = 0, n221 = 0, n222 = 0, n226 = 0, n227 = 0, n228 = 0;
reg n229 = 0, n230 = 0, n231 = 0, n232 = 0, n233 = 0, n234 = 0, n235 = 0, n236 = 0, n237 = 0, n238 = 0;
reg n246 = 0, n247 = 0, n248 = 0, n249 = 0, n250 = 0, n251 = 0, n252 = 0, n253 = 0, n254 = 0, n255 = 0;
reg n256 = 0, n257 = 0, n258 = 0, n259 = 0, n261 = 0, n262 = 0, io_13_31_0 = 0, n264 = 0, n265 = 0, n266 = 0;
reg n267 = 0, n268 = 0, n269 = 0, n270 = 0, n271 = 0, n272 = 0, n273 = 0, n274 = 0;
assign n289 = 1;
assign n473 = 1;

assign n288 =  1'b0;
assign n384 =  1'b0;
assign n395 =  1'b0;
assign n472 =  1'b0;
assign n277 =  !n79;
assign n278 =  (n184 ? 1'b0 : (n185 ? 1'b0 : n147));
assign n279 =  (n12 ? n51 : 1'b0);
assign n280 =  (n138 ? (n184 ? 1'b0 : !n185) : 1'b0);
assign n281 =  n18;
assign n282 =  n166;
assign n283 =  !n186;
assign n284 =  !n32;
assign n285 =  n272;
assign n286 =  (n12 ? !n248 : 1'b0);
assign n290 =  !n237;
assign n291 =  (n12 ? !n87 : 1'b0);
assign n292 =  (n12 ? !n16 : 1'b0);
assign n293 =  (n102 ? n12 : 1'b0);
assign n294 =  n41;
assign n295 =  !n54;
assign n296 =  (n109 ? n12 : 1'b0);
assign n297 =  (n160 ? n12 : 1'b0);
assign n298 =  (n175 ? 1'b0 : n12);
assign n299 =  n89;
assign n300 =  !n250;
assign n301 =  !n133;
assign n302 =  (n12 ? n135 : 1'b0);
assign n303 =  (n12 ? n238 : 1'b0);
assign n304 =  (n194 ? (n159 ? n149 : !n149) : (n159 ? !n149 : n149));
assign n305 =  !n90;
assign n306 =  !n103;
assign n307 =  (n12 ? !n55 : 1'b0);
assign n308 =  !io_16_0_0;
assign n309 =  !n45;
assign n310 =  !n222;
assign n311 =  (n240 ? !n226 : n226);
assign n312 =  (n185 ? 1'b0 : (n184 ? 1'b0 : (n12 ? !n144 : 1'b0)));
assign n313 =  (n15 ? 1'b0 : n12);
assign n314 =  !n53;
assign n315 =  !n75;
assign n316 =  !n81;
assign n317 =  (n12 ? n215 : 1'b0);
assign n318 =  n106;
assign n319 =  (n113 ? 1'b0 : n12);
assign n320 =  !n136;
assign n321 =  (n210 ? n12 : 1'b0);
assign n322 =  (n167 ? 1'b0 : n12);
assign n323 =  n93;
assign n324 =  (n12 ? !n96 : 1'b0);
assign n325 =  (n68 ? 1'b0 : n12);
assign n326 =  !n134;
assign n327 =  (n190 ? (n179 ? n159 : !n159) : (n179 ? !n159 : n159));
assign n328 =  (n201 ? (n159 ? n156 : !n156) : (n159 ? !n156 : n156));
assign n329 =  n198;
assign n330 =  n37;
assign n331 =  (n12 ? n28 : 1'b0);
assign n332 =  n257;
assign n333 =  n274;
assign n334 =  n67;
assign n335 =  (n242 ? !n228 : n228);
assign n336 =  n9;
assign n337 =  (n12 ? !n39 : 1'b0);
assign n338 =  (n43 ? n12 : 1'b0);
assign n339 =  n57;
assign n340 =  (n258 ? 1'b0 : n12);
assign n341 =  (n123 ? 1'b0 : n12);
assign n342 =  (n159 ? !n208 : n208);
assign n343 =  !n262;
assign n344 =  (n76 ? 1'b0 : n12);
assign n345 =  !n108;
assign n346 =  !n78;
assign n347 =  !n163;
assign n348 =  (n203 ? (n181 ? n159 : !n159) : (n181 ? !n159 : n159));
assign n349 =  (n192 ? (n159 ? n112 : !n112) : (n159 ? !n112 : n112));
assign n350 =  !n26;
assign n351 =  io_17_0_0;
assign n352 =  (n12 ? n49 : 1'b0);
assign n353 =  (n104 ? n12 : 1'b0);
assign n354 =  (n205 ? (n180 ? (n195 ? n155 : 1'b0) : 1'b0) : 1'b0);
assign n355 =  (n12 ? n220 : 1'b1);
assign n356 =  !n171;
assign n357 =  (n12 ? !n13 : 1'b0);
assign n358 =  !n60;
assign n359 =  (n12 ? !n35 : 1'b0);
assign n360 =  n125;
assign n361 =  (n244 ? !n230 : n230);
assign n362 =  (n211 ? n12 : 1'b0);
assign n363 =  (n12 ? !n168 : 1'b0);
assign n364 =  (n111 ? 1'b0 : n12);
assign n365 =  n91;
assign n366 =  !n94;
assign n367 =  (n185 ? 1'b0 : (n143 ? !n184 : 1'b0));
assign n368 =  n21;
assign n369 =  (n185 ? (n12 ? !n184 : 1'b1) : !n12);
assign n370 =  (n184 ? 1'b0 : (n185 ? 1'b0 : (n12 ? !n146 : 1'b0)));
assign n371 =  n70;
assign n372 =  n115;
assign n373 =  (n19 ? 1'b0 : n12);
assign n374 =  n66;
assign n375 =  !n31;
assign n376 =  (n40 ? 1'b0 : n12);
assign n377 =  !n266;
assign n378 =  (n12 ? !n110 : 1'b0);
assign n379 =  !n95;
assign n380 =  n249;
assign n381 =  (n12 ? !n107 : 1'b0);
assign n382 =  n82;
assign n385 =  !n119;
assign n386 =  (n12 ? !n56 : 1'b0);
assign n387 =  n232;
assign n388 =  (n12 ? n170 : 1'b0);
assign n389 =  !n216;
assign n390 =  !n153;
assign n391 =  !n50;
assign n392 =  !n151;
assign n393 =  n131;
assign n396 =  (n23 ? 1'b0 : n12);
assign n397 =  (n17 ? 1'b0 : n12);
assign n398 =  n36;
assign n399 =  n58;
assign n400 =  (n42 ? n12 : 1'b0);
assign n401 =  (n225 ? n223 : 1'b0);
assign n402 =  (n267 ? n12 : 1'b0);
assign n403 =  (n12 ? !n265 : 1'b0);
assign n404 =  !n271;
assign n405 =  (n141 ? 1'b0 : (n184 ? 1'b0 : (n185 ? 1'b0 : n12)));
assign n406 =  (n77 ? 1'b0 : n12);
assign n407 =  (n12 ? n218 : 1'b0);
assign n408 =  n65;
assign n409 =  (n92 ? 1'b0 : n12);
assign n410 =  n247;
assign n411 =  (n129 ? 1'b0 : n12);
assign n412 =  n83;
assign n413 =  (n189 ? (n150 ? n159 : !n159) : (n150 ? !n159 : n159));
assign n414 =  (n200 ? (n159 ? n158 : !n158) : (n159 ? !n158 : n158));
assign n415 =  !n268;
assign n416 =  (n52 ? n12 : 1'b0);
assign n417 =  (n12 ? (n184 ? 1'b1 : !n178) : 1'b1);
assign n418 =  (n105 ? n12 : 1'b0);
assign n419 =  (n183 ? (n184 ? 1'b0 : !n185) : 1'b0);
assign n420 =  n14;
assign n421 =  (n12 ? !n253 : 1'b0);
assign n422 =  (n184 ? 1'b0 : (n148 ? 1'b0 : (n12 ? !n185 : 1'b0)));
assign n423 =  n73;
assign n424 =  !n120;
assign n425 =  !n6;
assign n426 =  (n5 ? n12 : 1'b0);
assign n427 =  (n230 ? 1'b0 : (n208 ? 1'b0 : (n227 ? 1'b0 : !n222)));
assign n428 =  !n157;
assign n429 =  (n173 ? n12 : 1'b0);
assign n430 =  (n209 ? n12 : 1'b0);
assign n431 =  (n12 ? n213 : 1'b0);
assign n432 =  n71;
assign n433 =  (n84 ? 1'b0 : n12);
assign n434 =  (n12 ? !n130 : 1'b0);
assign n435 =  !n118;
assign n436 =  (n191 ? (n187 ? n159 : !n159) : (n187 ? !n159 : n159));
assign n437 =  n256;
assign n438 =  !n212;
assign n439 =  (n12 ? n236 : 1'b0);
assign n440 =  (n182 ? 1'b0 : (n177 ? 1'b0 : (n178 ? 1'b0 : n186)));
assign n441 =  (n255 ? 1'b0 : n12);
assign n442 =  n169;
assign n443 =  1'b1;
assign n444 =  n100;
assign n445 =  (n198 ? !io_16_0_0 : io_16_0_0);
assign n446 =  !n85;
assign n447 =  n124;
assign n448 =  n34;
assign n449 =  (n69 ? 1'b0 : n12);
assign n450 =  (n12 ? !n259 : 1'b0);
assign n451 =  (n101 ? n12 : 1'b0);
assign n452 =  (n234 ? 1'b0 : n12);
assign n453 =  !n154;
assign n454 =  (n161 ? n12 : 1'b0);
assign n455 =  (n12 ? !n174 : 1'b0);
assign n456 =  n22;
assign n457 =  (n127 ? 1'b0 : n12);
assign n458 =  (n193 ? (n159 ? n114 : !n114) : (n159 ? !n114 : n114));
assign n459 =  (n128 ? 1'b0 : n12);
assign n460 =  (n184 ? 1'b0 : (n185 ? 1'b0 : n137));
assign n461 =  (n149 ? 1'b0 : (n179 ? 1'b0 : (n181 ? 1'b0 : !n150)));
assign n462 =  !n219;
assign n463 =  !n8;
assign n464 =  !n152;
assign n465 =  !n132;
assign n466 =  (n264 ? 1'b0 : n12);
assign n467 =  (n184 ? 1'b0 : (n140 ? 1'b0 : (n12 ? !n185 : 1'b0)));
assign n468 =  n63;
assign n469 =  !n224;
assign n470 =  (n12 ? n122 : 1'b0);
assign n474 =  !n254;
assign n475 =  (n64 ? 1'b0 : n12);
assign n476 =  !n29;
assign n477 =  (n177 ? 1'b0 : (n185 ? 1'b0 : !n184));
assign n478 =  (n178 ? !n159 : n159);
assign n479 =  !n206;
assign n480 =  n74;
assign n481 =  !n121;
assign n482 =  (n11 ? 1'b0 : n12);
assign n483 =  (n46 ? n12 : 1'b0);
assign n484 =  (n228 ? (n231 ? (n226 ? n229 : 1'b0) : 1'b0) : 1'b0);
assign n485 =  (n12 ? n269 : 1'b0);
assign n486 =  (n241 ? !n227 : n227);
assign n487 =  (n12 ? (n185 ? 1'b0 : (n184 ? 1'b0 : !n142)) : 1'b0);
assign n488 =  (n12 ? n117 : 1'b0);
assign n489 =  (n12 ? !n273 : 1'b0);
assign n490 =  !n27;
assign n491 =  n88;
assign n492 =  n59;
assign n493 =  (n164 ? 1'b0 : n12);
assign n494 =  (n188 ? (n182 ? n159 : !n159) : (n182 ? !n159 : n159));
assign n495 =  n97;
assign n496 =  (n202 ? (n159 ? n197 : !n197) : (n159 ? !n197 : n197));
assign n497 =  !n217;
assign n498 =  !n7;
assign n499 =  n159;
assign n500 =  !n30;
assign n501 =  (n48 ? n12 : 1'b0);
assign n502 =  !n86;
assign n503 =  (n61 ? 1'b0 : n12);
assign n504 =  (n206 ? n153 : 1'b0);
assign n505 =  n126;
assign n506 =  !n251;
assign n507 =  (n270 ? n12 : 1'b0);
assign n508 =  (n98 ? 1'b0 : n12);
assign n509 =  (n157 ? (n152 ? (n151 ? n154 : 1'b0) : 1'b0) : 1'b0);
assign n510 =  (n243 ? !n229 : n229);
assign n511 =  !io_13_31_0;
assign n512 =  (n12 ? n261 : 1'b0);
assign n513 =  n33;
assign n514 =  (n25 ? n12 : 1'b0);
assign n515 =  n38;
assign n516 =  (n12 ? n116 : 1'b0);
assign n517 =  (n12 ? n80 : 1'b0);
assign n518 =  !n12;
assign n519 =  (n12 ? n235 : 1'b0);
assign n520 =  !n162;
assign n521 =  (n139 ? (n184 ? 1'b0 : !n185) : 1'b0);
assign n522 =  (n204 ? (n159 ? n199 : !n199) : (n159 ? !n199 : n199));
assign n523 =  !n172;
assign n524 =  n20;
assign n525 =  (n12 ? n47 : 1'b0);
assign n526 =  (n4 ? n12 : 1'b0);
assign n527 =  (n12 ? n252 : 1'b0);
assign n528 =  (n12 ? !n72 : 1'b0);
assign n529 =  (n245 ? !n231 : n231);
assign n530 =  n24;
assign n531 =  (n12 ? (n185 ? 1'b0 : (n184 ? 1'b0 : !n145)) : 1'b0);
assign n532 =  n10;
assign n533 =  (n12 ? n214 : 1'b0);
assign n534 =  (n165 ? 1'b0 : n12);
assign n535 =  (n12 ? n44 : 1'b0);
assign n536 =  n62;
assign n537 =  (n12 ? !n99 : 1'b0);
assign n538 =  (n233 ? 1'b0 : n12);
assign n539 =  (n198 ? !n221 : 1'b0);
assign n540 =  n246;
assign n275 =  (1'b0 & n208) | ((1'b0 | n208) & n289);
assign n200 =  (n149 & n159) | ((n149 | n159) & n194);
assign n241 =  (n226 & 1'b0) | ((n226 | 1'b0) & n240);
assign n191 =  (n159 & n179) | ((n159 | n179) & n190);
assign n202 =  (n156 & n159) | ((n156 | n159) & n201);
assign n243 =  (1'b0 & n228) | ((1'b0 | n228) & n242);
assign n204 =  (n159 & n181) | ((n159 | n181) & n203);
assign n193 =  (n112 & n159) | ((n112 | n159) & n192);
assign n245 =  (n230 & 1'b0) | ((n230 | 1'b0) & n244);
assign n188 =  (n177 & n159) | ((n177 | n159) & n276);
assign n240 =  (1'b0 & n222) | ((1'b0 | n222) & n275);
assign n190 =  (n159 & n150) | ((n159 | n150) & n189);
assign n201 =  (n158 & n159) | ((n158 | n159) & n200);
assign n192 =  (n159 & n187) | ((n159 | n187) & n191);
assign n194 =  (n114 & n159) | ((n114 | n159) & n193);
assign n276 =  (1'b0 & n178) | ((1'b0 | n178) & n473);
assign n242 =  (1'b0 & n227) | ((1'b0 | n227) & n241);
assign n189 =  (n159 & n182) | ((n159 | n182) & n188);
assign n203 =  (n197 & n159) | ((n197 | n159) & n202);
assign n244 =  (1'b0 & n229) | ((1'b0 | n229) & n243);
 always @(posedge io_12_31_1) if (n2) n82 <= n1 ? 1'b0 : n277;
 always @(posedge io_12_31_1) if (1'b1) n181 <= n1 ? 1'b0 : n278;
 always @(posedge io_12_31_1) if (n2) n47 <= n279;
 always @(posedge io_12_31_1) if (1'b1) n150 <= n1 ? 1'b0 : n280;
 always @(posedge io_12_31_1) if (n2) n17 <= n1 ? 1'b0 : n281;
 always @(posedge io_12_31_1) if (n2) n168 <= n1 ? 1'b0 : n282;
 assign n197 = n283;
 always @(posedge io_12_31_1) if (n2) n34 <= n1 ? 1'b0 : n284;
 always @(posedge io_12_31_1) if (n2) n274 <= n1 ? 1'b0 : n285;
 always @(posedge io_12_31_1) if (n2) n251 <= n286;
 assign n287 = n288;
 always @(posedge io_12_31_1) if (n2) n253 <= n1 ? 1'b0 : n290;
 always @(posedge io_12_31_1) if (n2) n85 <= n291;
 always @(posedge io_12_31_1) if (n2) n30 <= n292;
 always @(posedge io_12_31_1) if (n2) n103 <= n293;
 always @(posedge io_12_31_1) if (n2) n40 <= n1 ? 1'b0 : n294;
 always @(posedge io_12_31_1) if (n2) n55 <= n1 ? 1'b0 : n295;
 always @(posedge io_12_31_1) if (n2) n108 <= n296;
 always @(posedge io_12_31_1) if (n2) n163 <= n297;
 always @(posedge io_12_31_1) if (n2) n173 <= n298;
 always @(posedge io_12_31_1) if (n2) n106 <= n1 ? 1'b0 : n299;
 always @(posedge io_12_31_1) if (n2) n232 <= n1 ? 1'b0 : n300;
 always @(posedge io_12_31_1) if (n2) n128 <= n1 ? 1'b0 : n301;
 always @(posedge io_12_31_1) if (n2) n136 <= n302;
 always @(posedge io_12_31_1) if (n2) n254 <= n303;
 assign n143 = n304;
 always @(posedge io_12_31_1) if (n2) n87 <= n1 ? 1'b0 : n305;
 always @(posedge io_12_31_1) if (n2) n100 <= n1 ? 1'b0 : n306;
 always @(posedge io_12_31_1) if (n2) n49 <= n307;
 always @(posedge io_12_31_1) if (n196) n198 <= n1 ? 1'b0 : n308;
 always @(posedge io_12_31_1) if (n2) n68 <= n1 ? 1'b0 : n309;
 always @(posedge io_12_31_1) if (n208) n222 <= n310;
 always @(posedge io_12_31_1) if (n239) n226 <= n311;
 always @(posedge io_12_31_1) if (1'b1) n154 <= n312;
 always @(posedge io_12_31_1) if (n2) n32 <= n313;
 always @(posedge io_12_31_1) if (n2) n56 <= n1 ? 1'b0 : n314;
 always @(posedge io_12_31_1) if (n2) n57 <= n1 ? 1'b0 : n315;
 always @(posedge io_12_31_1) if (n2) n62 <= n1 ? 1'b0 : n316;
 always @(posedge io_12_31_1) if (n2) n219 <= n317;
 always @(posedge io_12_31_1) if (n2) n107 <= n1 ? 1'b0 : n318;
 always @(posedge io_12_31_1) if (n2) n117 <= n319;
 always @(posedge io_12_31_1) if (n2) n110 <= n1 ? 1'b0 : n320;
 always @(posedge io_12_31_1) if (n2) n212 <= n321;
 always @(posedge io_12_31_1) if (n2) n217 <= n322;
 always @(posedge io_12_31_1) if (n2) n77 <= n1 ? 1'b0 : n323;
 always @(posedge io_12_31_1) if (n2) n95 <= n324;
 always @(posedge io_12_31_1) if (n2) n81 <= n325;
 always @(posedge io_12_31_1) if (n2) n129 <= n1 ? 1'b0 : n326;
 assign n139 = n327;
 assign n145 = n328;
 always @(posedge io_12_31_1) if (1'b1) n221 <= n1 ? 1'b0 : n329;
 always @(posedge io_12_31_1) if (n2) n19 <= n1 ? 1'b0 : n330;
 always @(posedge io_12_31_1) if (n2) n51 <= n331;
 always @(posedge io_12_31_1) if (n2) n255 <= n1 ? 1'b0 : n332;
 always @(posedge io_12_31_1) if (n2) n273 <= n1 ? 1'b0 : n333;
 always @(posedge io_12_31_1) if (n2) n69 <= n1 ? 1'b0 : n334;
 always @(posedge io_12_31_1) if (n239) n228 <= n335;
 always @(posedge io_12_31_1) if (n2) n10 <= n1 ? 1'b0 : n336;
 always @(posedge io_12_31_1) if (n2) n25 <= n337;
 always @(posedge io_12_31_1) if (n2) n45 <= n338;
 always @(posedge io_12_31_1) if (n2) n59 <= n1 ? 1'b0 : n339;
 always @(posedge io_12_31_1) if (n2) n269 <= n340;
 always @(posedge io_12_31_1) if (n2) n118 <= n341;
 always @(posedge io_12_31_1) if (n239) n208 <= n342;
 always @(posedge io_12_31_1) if (n2) n246 <= n1 ? 1'b0 : n343;
 always @(posedge io_12_31_1) if (n2) n78 <= n344;
 always @(posedge io_12_31_1) if (n2) n92 <= n1 ? 1'b0 : n345;
 always @(posedge io_12_31_1) if (n2) n96 <= n1 ? 1'b0 : n346;
 always @(posedge io_12_31_1) if (n2) n130 <= n1 ? 1'b0 : n347;
 assign n147 = n348;
 assign n141 = n349;
 always @(posedge io_12_31_1) if (n2) n13 <= n1 ? 1'b0 : n350;
 always @(posedge io_12_31_1) if (n2) n259 <= n1 ? 1'b0 : n351;
 always @(posedge io_12_31_1) if (n2) n53 <= n352;
 always @(posedge io_12_31_1) if (n2) n90 <= n353;
 assign n185 = n354;
 assign n2 = n355;
 always @(posedge io_12_31_1) if (n2) n174 <= n1 ? 1'b0 : n356;
 always @(posedge io_12_31_1) if (n2) n28 <= n357;
 always @(posedge io_12_31_1) if (n2) n76 <= n1 ? 1'b0 : n358;
 always @(posedge io_12_31_1) if (n2) n29 <= n359;
 always @(posedge io_12_31_1) if (n2) n127 <= n1 ? 1'b0 : n360;
 always @(posedge io_12_31_1) if (n239) n230 <= n361;
 always @(posedge io_12_31_1) if (n2) n210 <= n362;
 always @(posedge io_12_31_1) if (n2) n214 <= n363;
 always @(posedge io_12_31_1) if (n2) n135 <= n364;
 always @(posedge io_12_31_1) if (n2) n93 <= n1 ? 1'b0 : n365;
 always @(posedge io_12_31_1) if (n2) n97 <= n1 ? 1'b0 : n366;
 always @(posedge io_12_31_1) if (1'b1) n149 <= n1 ? 1'b0 : n367;
 always @(posedge io_12_31_1) if (n2) n22 <= n1 ? 1'b0 : n368;
 assign n196 = n369;
 always @(posedge io_12_31_1) if (1'b1) n186 <= n370;
 always @(posedge io_12_31_1) if (n2) n67 <= n1 ? 1'b0 : n371;
 always @(posedge io_12_31_1) if (n2) n113 <= n1 ? 1'b0 : n372;
 always @(posedge io_12_31_1) if (n2) n4 <= n373;
 always @(posedge io_12_31_1) if (n2) n39 <= n1 ? 1'b0 : n374;
 always @(posedge io_12_31_1) if (n2) n35 <= n1 ? 1'b0 : n375;
 always @(posedge io_12_31_1) if (n2) n42 <= n376;
 always @(posedge io_12_31_1) if (n2) n265 <= n1 ? 1'b0 : n377;
 always @(posedge io_12_31_1) if (n2) n109 <= n378;
 always @(posedge io_12_31_1) if (n2) n91 <= n1 ? 1'b0 : n379;
 always @(posedge io_12_31_1) if (n2) n248 <= n1 ? 1'b0 : n380;
 always @(posedge io_12_31_1) if (n2) n132 <= n381;
 always @(posedge io_12_31_1) if (n2) n83 <= n1 ? 1'b0 : n382;
 assign n383 = n384;
 always @(posedge io_12_31_1) if (n2) n99 <= n1 ? 1'b0 : n385;
 always @(posedge io_12_31_1) if (n2) n48 <= n386;
 always @(posedge io_12_31_1) if (n2) n233 <= n1 ? 1'b0 : n387;
 always @(posedge io_12_31_1) if (n2) n235 <= n388;
 always @(posedge io_12_31_1) if (n2) n164 <= n1 ? 1'b0 : n389;
 assign n187 = n390;
 always @(posedge io_12_31_1) if (n2) n73 <= n1 ? 1'b0 : n391;
 assign n114 = n392;
 always @(posedge io_12_31_1) if (n2) n124 <= n1 ? 1'b0 : n393;
 assign n394 = n395;
 always @(posedge io_12_31_1) if (n2) n6 <= n396;
 always @(posedge io_12_31_1) if (n2) n31 <= n397;
 always @(posedge io_12_31_1) if (n2) n41 <= n1 ? 1'b0 : n398;
 always @(posedge io_12_31_1) if (n2) n36 <= n1 ? 1'b0 : n399;
 always @(posedge io_12_31_1) if (n2) n44 <= n400;
 assign n224 = n401;
 always @(posedge io_12_31_1) if (n2) n271 <= n402;
 always @(posedge io_12_31_1) if (n2) n267 <= n403;
 always @(posedge io_12_31_1) if (n2) n272 <= n1 ? 1'b0 : n404;
 always @(posedge io_12_31_1) if (1'b1) n152 <= n405;
 always @(posedge io_12_31_1) if (n2) n75 <= n406;
 always @(posedge io_12_31_1) if (n2) n216 <= n407;
 always @(posedge io_12_31_1) if (n2) n63 <= n1 ? 1'b0 : n408;
 always @(posedge io_12_31_1) if (n2) n94 <= n409;
 always @(posedge io_12_31_1) if (n2) n249 <= n1 ? 1'b0 : n410;
 always @(posedge io_12_31_1) if (n2) n133 <= n411;
 always @(posedge io_12_31_1) if (n2) n84 <= n1 ? 1'b0 : n412;
 assign n138 = n413;
 assign n144 = n414;
 always @(posedge io_12_31_1) if (n2) n257 <= n1 ? 1'b0 : n415;
 always @(posedge io_12_31_1) if (n2) n50 <= n416;
 assign n176 = n417;
 always @(posedge io_12_31_1) if (n2) n104 <= n418;
 always @(posedge io_12_31_1) if (1'b1) n178 <= n1 ? 1'b0 : n419;
 always @(posedge io_12_31_1) if (n2) n16 <= n1 ? 1'b0 : n420;
 always @(posedge io_12_31_1) if (n2) io_13_31_0 <= n421;
 always @(posedge io_12_31_1) if (1'b1) n206 <= n422;
 always @(posedge io_12_31_1) if (n2) n74 <= n1 ? 1'b0 : n423;
 always @(posedge io_12_31_1) if (n2) n115 <= n1 ? 1'b0 : n424;
 always @(posedge io_12_31_1) if (n2) n9 <= n1 ? 1'b0 : n425;
 always @(posedge io_12_31_1) if (n2) n7 <= n426;
 assign n225 = n427;
 assign n156 = n428;
 always @(posedge io_12_31_1) if (n2) n170 <= n429;
 always @(posedge io_12_31_1) if (n2) n213 <= n430;
 always @(posedge io_12_31_1) if (n2) n218 <= n431;
 always @(posedge io_12_31_1) if (n2) n65 <= n1 ? 1'b0 : n432;
 always @(posedge io_12_31_1) if (n2) n120 <= n433;
 always @(posedge io_12_31_1) if (n2) n134 <= n434;
 always @(posedge io_12_31_1) if (n2) n98 <= n1 ? 1'b0 : n435;
 assign n140 = n436;
 always @(posedge io_12_31_1) if (n2) n258 <= n1 ? 1'b0 : n437;
 always @(posedge io_12_31_1) if (n2) n234 <= n1 ? 1'b0 : n438;
 always @(posedge io_12_31_1) if (n2) n237 <= n439;
 assign n180 = n440;
 always @(posedge io_12_31_1) if (n2) n238 <= n441;
 always @(posedge io_12_31_1) if (n2) n167 <= n1 ? 1'b0 : n442;
 assign n159 = n443;
 always @(posedge io_12_31_1) if (n2) n111 <= n1 ? 1'b0 : n444;
 assign n184 = n445;
 always @(posedge io_12_31_1) if (n2) n70 <= n1 ? 1'b0 : n446;
 always @(posedge io_12_31_1) if (n2) n126 <= n1 ? 1'b0 : n447;
 always @(posedge io_12_31_1) if (n2) n33 <= n1 ? 1'b0 : n448;
 always @(posedge io_12_31_1) if (n2) n46 <= n449;
 always @(posedge io_12_31_1) if (n2) n270 <= n450;
 always @(posedge io_12_31_1) if (n2) n102 <= n451;
 always @(posedge io_12_31_1) if (n2) n209 <= n452;
 assign n158 = n453;
 always @(posedge io_12_31_1) if (n2) n162 <= n454;
 always @(posedge io_12_31_1) if (n2) n172 <= n455;
 always @(posedge io_12_31_1) if (n2) n24 <= n1 ? 1'b0 : n456;
 always @(posedge io_12_31_1) if (n2) n122 <= n457;
 assign n142 = n458;
 always @(posedge io_12_31_1) if (n2) n105 <= n459;
 always @(posedge io_12_31_1) if (1'b1) n182 <= n1 ? 1'b0 : n460;
 assign n195 = n461;
 always @(posedge io_12_31_1) if (n2) n169 <= n1 ? 1'b0 : n462;
 always @(posedge io_12_31_1) if (n2) n18 <= n1 ? 1'b0 : n463;
 assign n112 = n464;
 always @(posedge io_12_31_1) if (n2) n175 <= n1 ? 1'b0 : n465;
 always @(posedge io_12_31_1) if (n2) n252 <= n466;
 always @(posedge io_12_31_1) if (1'b1) n153 <= n467;
 always @(posedge io_12_31_1) if (n2) n61 <= n1 ? 1'b0 : n468;
 assign n239 = n469;
 always @(posedge io_12_31_1) if (n2) n116 <= n470;
 assign n471 = n472;
 always @(posedge io_12_31_1) if (n2) n256 <= n1 ? 1'b0 : n474;
 always @(posedge io_12_31_1) if (n2) n80 <= n475;
 always @(posedge io_12_31_1) if (n2) n14 <= n1 ? 1'b0 : n476;
 always @(posedge io_12_31_1) if (n176) n177 <= n1 ? 1'b0 : n477;
 assign n183 = n478;
 assign n199 = n479;
 always @(posedge io_12_31_1) if (n2) n72 <= n1 ? 1'b0 : n480;
 always @(posedge io_12_31_1) if (n2) n123 <= n1 ? 1'b0 : n481;
 always @(posedge io_12_31_1) if (n2) n5 <= n482;
 always @(posedge io_12_31_1) if (n2) n43 <= n483;
 assign n223 = n484;
 always @(posedge io_12_31_1) if (n2) n266 <= n485;
 always @(posedge io_12_31_1) if (n239) n227 <= n486;
 always @(posedge io_12_31_1) if (1'b1) n151 <= n487;
 always @(posedge io_12_31_1) if (n2) n160 <= n488;
 always @(posedge io_12_31_1) if (n2) n261 <= n489;
 always @(posedge io_12_31_1) if (n2) n23 <= n1 ? 1'b0 : n490;
 always @(posedge io_12_31_1) if (n2) n89 <= n1 ? 1'b0 : n491;
 always @(posedge io_12_31_1) if (n2) n58 <= n1 ? 1'b0 : n492;
 always @(posedge io_12_31_1) if (n2) n215 <= n493;
 assign n137 = n494;
 always @(posedge io_12_31_1) if (n2) n71 <= n1 ? 1'b0 : n495;
 assign n146 = n496;
 always @(posedge io_12_31_1) if (n2) n165 <= n1 ? 1'b0 : n497;
 always @(posedge io_12_31_1) if (n2) n15 <= n1 ? 1'b0 : n498;
 always @(posedge io_12_31_1) if (n224) n12 <= n499;
 always @(posedge io_12_31_1) if (n2) n20 <= n1 ? 1'b0 : n500;
 always @(posedge io_12_31_1) if (n2) n52 <= n501;
 always @(posedge io_12_31_1) if (n2) n88 <= n1 ? 1'b0 : n502;
 always @(posedge io_12_31_1) if (n2) n60 <= n503;
 assign n205 = n504;
 always @(posedge io_12_31_1) if (n2) n125 <= n1 ? 1'b0 : n505;
 always @(posedge io_12_31_1) if (n2) n264 <= n1 ? 1'b0 : n506;
 always @(posedge io_12_31_1) if (n2) n268 <= n507;
 always @(posedge io_12_31_1) if (n2) n101 <= n508;
 assign n155 = n509;
 always @(posedge io_12_31_1) if (n239) n229 <= n510;
 assign io_17_0_0 = n511;
 always @(posedge io_12_31_1) if (n2) n262 <= n512;
 always @(posedge io_12_31_1) if (n2) n37 <= n1 ? 1'b0 : n513;
 always @(posedge io_12_31_1) if (n2) n26 <= n514;
 always @(posedge io_12_31_1) if (n2) n64 <= n1 ? 1'b0 : n515;
 always @(posedge io_12_31_1) if (n2) n119 <= n516;
 always @(posedge io_12_31_1) if (n2) n79 <= n517;
 assign n1 = n518;
 always @(posedge io_12_31_1) if (n2) n236 <= n519;
 always @(posedge io_12_31_1) if (n2) n131 <= n1 ? 1'b0 : n520;
 always @(posedge io_12_31_1) if (1'b1) n179 <= n1 ? 1'b0 : n521;
 assign n148 = n522;
 always @(posedge io_12_31_1) if (n2) n166 <= n1 ? 1'b0 : n523;
 always @(posedge io_12_31_1) if (n2) n21 <= n1 ? 1'b0 : n524;
 always @(posedge io_12_31_1) if (n2) n54 <= n525;
 always @(posedge io_12_31_1) if (n2) n8 <= n526;
 always @(posedge io_12_31_1) if (n2) n250 <= n527;
 always @(posedge io_12_31_1) if (n2) n86 <= n528;
 always @(posedge io_12_31_1) if (n239) n231 <= n529;
 always @(posedge io_12_31_1) if (n2) n38 <= n1 ? 1'b0 : n530;
 always @(posedge io_12_31_1) if (1'b1) n157 <= n531;
 always @(posedge io_12_31_1) if (n2) n11 <= n1 ? 1'b0 : n532;
 always @(posedge io_12_31_1) if (n2) n161 <= n533;
 always @(posedge io_12_31_1) if (n2) n171 <= n534;
 always @(posedge io_12_31_1) if (n2) n27 <= n535;
 always @(posedge io_12_31_1) if (n2) n66 <= n1 ? 1'b0 : n536;
 always @(posedge io_12_31_1) if (n2) n121 <= n537;
 always @(posedge io_12_31_1) if (n2) n211 <= n538;
 always @(posedge io_12_31_1) if (1'b1) n220 <= n1 ? 1'b0 : n539;
 always @(posedge io_12_31_1) if (n2) n247 <= n1 ? 1'b0 : n540;

endmodule

